------------------------- 1. 2x1 mux ----------------------------------
library ieee;
USE ieee.std_logic_1164.all;
-----------------------------------------------------------------------
ENTITY mux is
    PORT(
        a,b,sel : IN std_logic;
        y : OUT std_logic
    );
-----------------------------------------------------------------------
architecture mux OF mux is
begin
    when (sel = '0') => y = a;
    when (sel = '1') => y = b;
end mux;

--- 3. 7segment decoder 
--- 4. mux를 활용해 5개의 3비트를 제공. 이들 중 하나를 mux를 활용해 출력해라.


--- 1. 2진수를  10진수로 변환해라.(10 이상 포함) if, else 구문 활용 
--- 1. 2진수를  10진수로 변환해라.(10 이상 포함) if, else 구문 활용 X
--- 2. 가산기 제작
--- 3. 4bit 가산기 제작
--- 5. 4bit 2진수 2개를 더해 10진수로 표현하라
